module KeyGenerator(
    input [127:0] Key,
    input fOdd,
    output [63:0] o_Key
);



endmodule