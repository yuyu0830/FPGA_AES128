module UART_Top()